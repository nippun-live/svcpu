`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/03/2024 07:09:00 PM
// Design Name: 
// Module Name: databus_mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module databus_mux( input logic [15:0] din_MARMUX, din_PC, din_ALU, din_MDR, 
                    input logic [1:0] select, 
                    output logic [15:0] dout );
                    
always_comb
begin
dout = 16'b0;
if (select == 2'b00) 
    begin
    dout = din_MARMUX; 
    end
else if (select == 2'b01)
    begin
    dout = din_PC;
    end
else if (select == 2'b10)
    begin
    dout = din_ALU;
    end
else if (select == 2'b11)
    begin
    dout = din_MDR;
    end
else
    begin
    dout = 16'b0;
    end

end
endmodule